library verilog;
use verilog.vl_types.all;
entity bilinear_vlg_tst is
end bilinear_vlg_tst;
